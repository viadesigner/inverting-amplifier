
* Project OPAMP
* Mentor Graphics Netlist Created with Version 5.8
* File created Mon Feb 25 11:25:06 2013
* Inifile   : 
*
* Config file: C:\MentorGraphics\SystemVision5.9\standard\svspice.cfg
*
* Options   : -_ -h -kC:\MentorGraphics\SystemVision5.9\standard\svspice.cfg -gopamp.tempfile 
* 
* Levels    : 
* 
.option noinclib
* Models for Eldo<->VHDL-AMS data conversion
.model a2d_eldo a2d mode=std_logic VTH=1.65
.model d2a_eldo d2a mode=std_logic VHI=3.3 VLO=0.0
.defhook a2d_eldo
.defhook d2a_eldo
.param process_corner=0
YAMP2 VIA_AMP_OA(LEVEL_2) GENERIC: AVOL="(102.3,92.9,100.1)" AVOL_NOM="102" 
+ CMRR="(104.8,96.0,104.3)" FPARA="(59.0,225.0,5.5)" FZC="(48.6,202.0,35.5)" 
+ FZP="(0.096,0.595,0.0846)" IBIAS="(10.0,18.45,6.1)" IDD_NOM="737" 
+ ISRATIO="(73.7,73.7,73.7)" PSRR="(98.0,87.5,94.0)" ROUT="(0.95,0.6,1.6)" 
+ SR="(23.3,42.9,13.1)" SR_NOM="23" TC_AVOL="(-1273,-1273,-1273)" 
+ TC_CMRR="(-807,-807,-807)" TC_FPARA="(-7954,-7954,-7954)" 
+ TC_FZC="(8042,8042,8042)" TC_FZP="(6286,6286,6286)" 
+ TC_PSRR="(-1496,-1496,-1496)" TC_ROUT="(3047,3047,3047)" 
+ TC_SR="(-1084,-1084,-1084)" TC_UGB="(-2982,-2982,-2982)" 
+ UGB="(11.7,26.0,6.33)" UGB_NOM="12" VOS_MAX="0.013" 
+ VOS_MISMATCH="(0.0133,0.0133,0.0133)" PORT: VCM N1N4 AVDD AVDD AVSS VOUT
YV1 V_CONSTANT(IDEAL) GENERIC: LEVEL="0.0" PORT: AVSS 0
YV_SINE1 V_SINE(IDEAL) GENERIC: AMPLITUDE="0.5" FREQ="500.0" PORT: VIN VCM
YV2 V_CONSTANT(IDEAL) GENERIC: LEVEL="1.65" PORT: VCM AVSS
YV3 V_CONSTANT(IDEAL) GENERIC: LEVEL="1.65" PORT: AVDD VCM
YR3 VIA_RES_2P(LEVEL_2) GENERIC: 
+ ACTUALRESISTANCE="(6500.0,5200.0,7913.04347826)" AREA="48" 
+ PARASITICA="(4.97E-15,4.05E-15,8.5E-15)" 
+ PARASITICA2ABOVE="(2.42E-15,1.68E-15,5.71E-15)" 
+ PARASITICA2BELOW="(2.55E-15,2.37E-15,2.79E-15)" 
+ PARASITICB="(4.97E-15,4.05E-15,8.5E-15)" 
+ PARASITICB2ABOVE="(2.42E-15,1.68E-15,5.71E-15)" 
+ PARASITICB2BELOW="(2.55E-15,2.37E-15,2.79E-15)" PORT: VIN N1N4
YR4 VIA_RES_2P(LEVEL_2) GENERIC: 
+ ACTUALRESISTANCE="(13000.0,10400.0,15826.0869565)" AREA="97" 
+ AREARESISTORTOTAL="67.6" DESIREDRESISTANCE="13E3" NOMINALRESISTANCE="13000" 
+ NUMUNITRESISTORS="2" PARASITICA="(9.94E-15,8.1E-15,1.7E-14)" 
+ PARASITICA2ABOVE="(4.84E-15,3.36E-15,1.142E-14)" 
+ PARASITICA2BELOW="(5.1E-15,4.74E-15,5.58E-15)" 
+ PARASITICB="(9.94E-15,8.1E-15,1.7E-14)" 
+ PARASITICB2ABOVE="(4.84E-15,3.36E-15,1.142E-14)" 
+ PARASITICB2BELOW="(5.1E-15,4.74E-15,5.58E-15)" PORT: N1N4 VOUT
* DICTIONARY 1
* GND = 0
.GLOBAL ELECTRICAL_REF
.model VIA_RES_2P(LEVEL_2) macro lang=vhdlams LIB=WORK
.model V_CONSTANT(IDEAL) macro lang=vhdlams LIB=EDULIB
.model VIA_AMP_OA(LEVEL_2) macro lang=vhdlams LIB=WORK
.model V_SINE(IDEAL) macro lang=vhdlams LIB=EDULIB
.END
